library verilog;
use verilog.vl_types.all;
entity tb_half_adder is
end tb_half_adder;
