library verilog;
use verilog.vl_types.all;
entity tb_state_machine is
end tb_state_machine;
