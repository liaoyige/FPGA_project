library verilog;
use verilog.vl_types.all;
entity tb_decoder is
end tb_decoder;
