library verilog;
use verilog.vl_types.all;
entity tb_flip_flop is
end tb_flip_flop;
