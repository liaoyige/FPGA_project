library verilog;
use verilog.vl_types.all;
entity tb_divider_six is
end tb_divider_six;
