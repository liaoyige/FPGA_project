library verilog;
use verilog.vl_types.all;
entity tb_full_adder_top is
end tb_full_adder_top;
