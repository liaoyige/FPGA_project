library verilog;
use verilog.vl_types.all;
entity tb_pll is
end tb_pll;
