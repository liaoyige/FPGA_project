library verilog;
use verilog.vl_types.all;
entity tb_state_machine_up_1 is
end tb_state_machine_up_1;
