library verilog;
use verilog.vl_types.all;
entity tb_divider_five is
end tb_divider_five;
